module simutest(c, a, b);
output c;
input a, b;

assign c = a&b;
endmodule 