module test(c, a, b);
output c;
input a, b;

    xor G1(c, a, b);
//    and G1(c, a, b);
endmodule
