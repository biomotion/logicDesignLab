module flipflop()
endmodule
